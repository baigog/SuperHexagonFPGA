library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY CONTROLADOR_VGA IS
	PORT(
		CLK		:	IN	STD_LOGIC;
		CLR		:	IN	STD_LOGIC;
		RED_IN	:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN_IN	:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE_IN	:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		
		HSYNC		:	OUT	STD_LOGIC;
		VSYNC		:	OUT	STD_LOGIC;
		X			:	OUT	UNSIGNED(9 DOWNTO 0);
		Y			:	OUT	UNSIGNED(9 DOWNTO 0);
		RED		:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN		:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE		:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		END_FRAME:	OUT	STD_LOGIC;
		PRE_FRAME:	OUT	STD_LOGIC
		);
END ENTITY;

ARCHITECTURE BEH OF CONTROLADOR_VGA IS

CONSTANT PX_DLY	: UNSIGNED:= TO_UNSIGNED(2,10);
CONSTANT HPIXELS	: UNSIGNED:= TO_UNSIGNED(800,10);
CONSTANT vLINES	: UNSIGNED:= TO_UNSIGNED(521,10);
CONSTANT HPULSE	: UNSIGNED:= TO_UNSIGNED(96,10);
CONSTANT VPULSE	: UNSIGNED:= TO_UNSIGNED(2,10);
CONSTANT HBP		: UNSIGNED:= TO_UNSIGNED(144,10);
CONSTANT HFP		: UNSIGNED:= TO_UNSIGNED(784,10);
CONSTANT VBP		: UNSIGNED:= TO_UNSIGNED(31,10);
CONSTANT VFP		: UNSIGNED:= TO_UNSIGNED(511,10);

SIGNAL	HC	:	UNSIGNED(9 DOWNTO 0);
SIGNAL	VC	:	UNSIGNED(9 DOWNTO 0);
SIGNAL	IN_FRAME	:	STD_LOGIC;

BEGIN

HSYNC<='0' WHEN (HC<HPULSE) ELSE '1';
VSYNC<='0' WHEN (VC<VPULSE) ELSE '1';
IN_FRAME <= '1' WHEN ((VC >= VBP AND VC < VFP) AND (HC >= HBP AND HC < (HBP+TO_UNSIGNED(640,10)))) ELSE '0';
PRE_FRAME <= '1' WHEN (HC=(9 DOWNTO 0 => '0') AND VC=(9 DOWNTO 0 => '0')) ELSE '0';
END_FRAME <= '1' WHEN (HC=(9 DOWNTO 0 => '0') AND VC=TO_UNSIGNED(515,10)) ELSE '0';

SUMACONTADORES:PROCESS (CLK,CLR,HC,VC)
BEGIN
IF (CLR='1') THEN
	HC<=(OTHERS=>'0');
	VC<=(OTHERS=>'0');
ELSIF (RISING_EDGE(CLK)) THEN
	IF(HC < HPIXELS-1) THEN
		HC<=HC+1;
	ELSE
		HC<=(OTHERS=>'0');
		IF(VC < VLINES-1) THEN
			VC<=VC+1;
		ELSE
			VC<=(OTHERS=>'0');
		END IF;
	END IF;
END IF;
END PROCESS;

SETEACOORDENADAS:PROCESS (CLK,VC,HC)
BEGIN
	IF(RISING_EDGE(CLK)) THEN
		IF(VC >= VBP AND VC < VFP) THEN
			Y <= VC-VBP;
		ELSE
			Y <= (OTHERS=>'0');
		END IF;
		IF(HC >= HBP - PX_DLY AND HC < (HBP+TO_UNSIGNED(640,10)-PX_DLY)) THEN
		X <= HC+PX_DLY-HBP;
		ELSE
			X	<=	(OTHERS=>'0');
		END IF;
	END IF;
END PROCESS;

SETEACOLORES:PROCESS (CLK,IN_FRAME)
BEGIN
IF RISING_EDGE(CLK) THEN
	IF (IN_FRAME='1') THEN
		RED <= RED_IN;
		GREEN <= GREEN_IN;
		BLUE <= BLUE_IN;
	ELSE
		RED <= (OTHERS => '0');
		GREEN <= (OTHERS => '0');
		BLUE <= (OTHERS => '0');
	END IF;
END IF;
END PROCESS;

END ARCHITECTURE;
