library ieee;
use ieee.std_logic_1164.all;

ENTITY PRUEBA_VGA IS
	PORT(
		CLK	:	IN		STD_LOGIC;
		X		:	IN		STD_LOGIC_VECTOR(9 DOWNTO 0);
		Y		:	IN		STD_LOGIC_VECTOR(9 DOWNTO 0);
		RED	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEH OF PRUEBA_VGA IS
BEGIN

PROCESS (CLK)
BEGIN
	IF (RISING_EDGE(CLK)) THEN
		RED <= X(4 DOWNTO 1);
		GREEN <= Y(4 DOWNTO 1);
		BLUE(1 DOWNTO 0) <= X(6 DOWNTO 5);
		BLUE(3 DOWNTO 2) <= X(6 DOWNTO 5);
	END IF;
END PROCESS;

END ARCHITECTURE;